library verilog;
use verilog.vl_types.all;
entity IC_8259A_DUT is
end IC_8259A_DUT;
